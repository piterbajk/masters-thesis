// multicore_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module multicore_system (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         core_0_data_master_waitrequest;                  // mm_interconnect_0:core_0_data_master_waitrequest -> core_0:data_master_waitrequest
	wire  [31:0] core_0_data_master_readdata;                     // mm_interconnect_0:core_0_data_master_readdata -> core_0:data_master_readdata
	wire         core_0_data_master_debugaccess;                  // core_0:data_master_debugaccess -> mm_interconnect_0:core_0_data_master_debugaccess
	wire  [19:0] core_0_data_master_address;                      // core_0:data_master_address -> mm_interconnect_0:core_0_data_master_address
	wire         core_0_data_master_read;                         // core_0:data_master_read -> mm_interconnect_0:core_0_data_master_read
	wire   [3:0] core_0_data_master_byteenable;                   // core_0:data_master_byteenable -> mm_interconnect_0:core_0_data_master_byteenable
	wire         core_0_data_master_readdatavalid;                // mm_interconnect_0:core_0_data_master_readdatavalid -> core_0:data_master_readdatavalid
	wire  [31:0] core_0_data_master_writedata;                    // core_0:data_master_writedata -> mm_interconnect_0:core_0_data_master_writedata
	wire         core_0_data_master_write;                        // core_0:data_master_write -> mm_interconnect_0:core_0_data_master_write
	wire   [0:0] core_0_data_master_burstcount;                   // core_0:data_master_burstcount -> mm_interconnect_0:core_0_data_master_burstcount
	wire         core_1_data_master_waitrequest;                  // mm_interconnect_0:core_1_data_master_waitrequest -> core_1:data_master_waitrequest
	wire  [31:0] core_1_data_master_readdata;                     // mm_interconnect_0:core_1_data_master_readdata -> core_1:data_master_readdata
	wire         core_1_data_master_debugaccess;                  // core_1:data_master_debugaccess -> mm_interconnect_0:core_1_data_master_debugaccess
	wire  [19:0] core_1_data_master_address;                      // core_1:data_master_address -> mm_interconnect_0:core_1_data_master_address
	wire         core_1_data_master_read;                         // core_1:data_master_read -> mm_interconnect_0:core_1_data_master_read
	wire   [3:0] core_1_data_master_byteenable;                   // core_1:data_master_byteenable -> mm_interconnect_0:core_1_data_master_byteenable
	wire         core_1_data_master_readdatavalid;                // mm_interconnect_0:core_1_data_master_readdatavalid -> core_1:data_master_readdatavalid
	wire  [31:0] core_1_data_master_writedata;                    // core_1:data_master_writedata -> mm_interconnect_0:core_1_data_master_writedata
	wire         core_1_data_master_write;                        // core_1:data_master_write -> mm_interconnect_0:core_1_data_master_write
	wire   [0:0] core_1_data_master_burstcount;                   // core_1:data_master_burstcount -> mm_interconnect_0:core_1_data_master_burstcount
	wire         core_2_data_master_waitrequest;                  // mm_interconnect_0:core_2_data_master_waitrequest -> core_2:data_master_waitrequest
	wire  [31:0] core_2_data_master_readdata;                     // mm_interconnect_0:core_2_data_master_readdata -> core_2:data_master_readdata
	wire         core_2_data_master_debugaccess;                  // core_2:data_master_debugaccess -> mm_interconnect_0:core_2_data_master_debugaccess
	wire  [19:0] core_2_data_master_address;                      // core_2:data_master_address -> mm_interconnect_0:core_2_data_master_address
	wire         core_2_data_master_read;                         // core_2:data_master_read -> mm_interconnect_0:core_2_data_master_read
	wire   [3:0] core_2_data_master_byteenable;                   // core_2:data_master_byteenable -> mm_interconnect_0:core_2_data_master_byteenable
	wire         core_2_data_master_readdatavalid;                // mm_interconnect_0:core_2_data_master_readdatavalid -> core_2:data_master_readdatavalid
	wire  [31:0] core_2_data_master_writedata;                    // core_2:data_master_writedata -> mm_interconnect_0:core_2_data_master_writedata
	wire         core_2_data_master_write;                        // core_2:data_master_write -> mm_interconnect_0:core_2_data_master_write
	wire   [0:0] core_2_data_master_burstcount;                   // core_2:data_master_burstcount -> mm_interconnect_0:core_2_data_master_burstcount
	wire         core_7_data_master_waitrequest;                  // mm_interconnect_0:core_7_data_master_waitrequest -> core_7:data_master_waitrequest
	wire  [31:0] core_7_data_master_readdata;                     // mm_interconnect_0:core_7_data_master_readdata -> core_7:data_master_readdata
	wire         core_7_data_master_debugaccess;                  // core_7:data_master_debugaccess -> mm_interconnect_0:core_7_data_master_debugaccess
	wire  [19:0] core_7_data_master_address;                      // core_7:data_master_address -> mm_interconnect_0:core_7_data_master_address
	wire         core_7_data_master_read;                         // core_7:data_master_read -> mm_interconnect_0:core_7_data_master_read
	wire   [3:0] core_7_data_master_byteenable;                   // core_7:data_master_byteenable -> mm_interconnect_0:core_7_data_master_byteenable
	wire         core_7_data_master_readdatavalid;                // mm_interconnect_0:core_7_data_master_readdatavalid -> core_7:data_master_readdatavalid
	wire  [31:0] core_7_data_master_writedata;                    // core_7:data_master_writedata -> mm_interconnect_0:core_7_data_master_writedata
	wire         core_7_data_master_write;                        // core_7:data_master_write -> mm_interconnect_0:core_7_data_master_write
	wire   [0:0] core_7_data_master_burstcount;                   // core_7:data_master_burstcount -> mm_interconnect_0:core_7_data_master_burstcount
	wire         core_3_data_master_waitrequest;                  // mm_interconnect_0:core_3_data_master_waitrequest -> core_3:data_master_waitrequest
	wire  [31:0] core_3_data_master_readdata;                     // mm_interconnect_0:core_3_data_master_readdata -> core_3:data_master_readdata
	wire         core_3_data_master_debugaccess;                  // core_3:data_master_debugaccess -> mm_interconnect_0:core_3_data_master_debugaccess
	wire  [19:0] core_3_data_master_address;                      // core_3:data_master_address -> mm_interconnect_0:core_3_data_master_address
	wire         core_3_data_master_read;                         // core_3:data_master_read -> mm_interconnect_0:core_3_data_master_read
	wire   [3:0] core_3_data_master_byteenable;                   // core_3:data_master_byteenable -> mm_interconnect_0:core_3_data_master_byteenable
	wire         core_3_data_master_readdatavalid;                // mm_interconnect_0:core_3_data_master_readdatavalid -> core_3:data_master_readdatavalid
	wire  [31:0] core_3_data_master_writedata;                    // core_3:data_master_writedata -> mm_interconnect_0:core_3_data_master_writedata
	wire         core_3_data_master_write;                        // core_3:data_master_write -> mm_interconnect_0:core_3_data_master_write
	wire   [0:0] core_3_data_master_burstcount;                   // core_3:data_master_burstcount -> mm_interconnect_0:core_3_data_master_burstcount
	wire         core_4_data_master_waitrequest;                  // mm_interconnect_0:core_4_data_master_waitrequest -> core_4:data_master_waitrequest
	wire  [31:0] core_4_data_master_readdata;                     // mm_interconnect_0:core_4_data_master_readdata -> core_4:data_master_readdata
	wire         core_4_data_master_debugaccess;                  // core_4:data_master_debugaccess -> mm_interconnect_0:core_4_data_master_debugaccess
	wire  [19:0] core_4_data_master_address;                      // core_4:data_master_address -> mm_interconnect_0:core_4_data_master_address
	wire         core_4_data_master_read;                         // core_4:data_master_read -> mm_interconnect_0:core_4_data_master_read
	wire   [3:0] core_4_data_master_byteenable;                   // core_4:data_master_byteenable -> mm_interconnect_0:core_4_data_master_byteenable
	wire         core_4_data_master_readdatavalid;                // mm_interconnect_0:core_4_data_master_readdatavalid -> core_4:data_master_readdatavalid
	wire  [31:0] core_4_data_master_writedata;                    // core_4:data_master_writedata -> mm_interconnect_0:core_4_data_master_writedata
	wire         core_4_data_master_write;                        // core_4:data_master_write -> mm_interconnect_0:core_4_data_master_write
	wire   [0:0] core_4_data_master_burstcount;                   // core_4:data_master_burstcount -> mm_interconnect_0:core_4_data_master_burstcount
	wire         core_5_data_master_waitrequest;                  // mm_interconnect_0:core_5_data_master_waitrequest -> core_5:data_master_waitrequest
	wire  [31:0] core_5_data_master_readdata;                     // mm_interconnect_0:core_5_data_master_readdata -> core_5:data_master_readdata
	wire         core_5_data_master_debugaccess;                  // core_5:data_master_debugaccess -> mm_interconnect_0:core_5_data_master_debugaccess
	wire  [19:0] core_5_data_master_address;                      // core_5:data_master_address -> mm_interconnect_0:core_5_data_master_address
	wire         core_5_data_master_read;                         // core_5:data_master_read -> mm_interconnect_0:core_5_data_master_read
	wire   [3:0] core_5_data_master_byteenable;                   // core_5:data_master_byteenable -> mm_interconnect_0:core_5_data_master_byteenable
	wire         core_5_data_master_readdatavalid;                // mm_interconnect_0:core_5_data_master_readdatavalid -> core_5:data_master_readdatavalid
	wire  [31:0] core_5_data_master_writedata;                    // core_5:data_master_writedata -> mm_interconnect_0:core_5_data_master_writedata
	wire         core_5_data_master_write;                        // core_5:data_master_write -> mm_interconnect_0:core_5_data_master_write
	wire   [0:0] core_5_data_master_burstcount;                   // core_5:data_master_burstcount -> mm_interconnect_0:core_5_data_master_burstcount
	wire         core_6_data_master_waitrequest;                  // mm_interconnect_0:core_6_data_master_waitrequest -> core_6:data_master_waitrequest
	wire  [31:0] core_6_data_master_readdata;                     // mm_interconnect_0:core_6_data_master_readdata -> core_6:data_master_readdata
	wire         core_6_data_master_debugaccess;                  // core_6:data_master_debugaccess -> mm_interconnect_0:core_6_data_master_debugaccess
	wire  [19:0] core_6_data_master_address;                      // core_6:data_master_address -> mm_interconnect_0:core_6_data_master_address
	wire         core_6_data_master_read;                         // core_6:data_master_read -> mm_interconnect_0:core_6_data_master_read
	wire   [3:0] core_6_data_master_byteenable;                   // core_6:data_master_byteenable -> mm_interconnect_0:core_6_data_master_byteenable
	wire         core_6_data_master_readdatavalid;                // mm_interconnect_0:core_6_data_master_readdatavalid -> core_6:data_master_readdatavalid
	wire  [31:0] core_6_data_master_writedata;                    // core_6:data_master_writedata -> mm_interconnect_0:core_6_data_master_writedata
	wire         core_6_data_master_write;                        // core_6:data_master_write -> mm_interconnect_0:core_6_data_master_write
	wire   [0:0] core_6_data_master_burstcount;                   // core_6:data_master_burstcount -> mm_interconnect_0:core_6_data_master_burstcount
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;  // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;   // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_core_1_mailbox_in_readdata;    // core_1:mailbox_in_readdata -> mm_interconnect_0:core_1_mailbox_in_readdata
	wire         mm_interconnect_0_core_1_mailbox_in_waitrequest; // core_1:mailbox_in_waitrequest -> mm_interconnect_0:core_1_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_1_mailbox_in_address;     // mm_interconnect_0:core_1_mailbox_in_address -> core_1:mailbox_in_address
	wire         mm_interconnect_0_core_1_mailbox_in_read;        // mm_interconnect_0:core_1_mailbox_in_read -> core_1:mailbox_in_read
	wire         mm_interconnect_0_core_1_mailbox_in_write;       // mm_interconnect_0:core_1_mailbox_in_write -> core_1:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_1_mailbox_in_writedata;   // mm_interconnect_0:core_1_mailbox_in_writedata -> core_1:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_2_mailbox_in_readdata;    // core_2:mailbox_in_readdata -> mm_interconnect_0:core_2_mailbox_in_readdata
	wire         mm_interconnect_0_core_2_mailbox_in_waitrequest; // core_2:mailbox_in_waitrequest -> mm_interconnect_0:core_2_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_2_mailbox_in_address;     // mm_interconnect_0:core_2_mailbox_in_address -> core_2:mailbox_in_address
	wire         mm_interconnect_0_core_2_mailbox_in_read;        // mm_interconnect_0:core_2_mailbox_in_read -> core_2:mailbox_in_read
	wire         mm_interconnect_0_core_2_mailbox_in_write;       // mm_interconnect_0:core_2_mailbox_in_write -> core_2:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_2_mailbox_in_writedata;   // mm_interconnect_0:core_2_mailbox_in_writedata -> core_2:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_3_mailbox_in_readdata;    // core_3:mailbox_in_readdata -> mm_interconnect_0:core_3_mailbox_in_readdata
	wire         mm_interconnect_0_core_3_mailbox_in_waitrequest; // core_3:mailbox_in_waitrequest -> mm_interconnect_0:core_3_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_3_mailbox_in_address;     // mm_interconnect_0:core_3_mailbox_in_address -> core_3:mailbox_in_address
	wire         mm_interconnect_0_core_3_mailbox_in_read;        // mm_interconnect_0:core_3_mailbox_in_read -> core_3:mailbox_in_read
	wire         mm_interconnect_0_core_3_mailbox_in_write;       // mm_interconnect_0:core_3_mailbox_in_write -> core_3:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_3_mailbox_in_writedata;   // mm_interconnect_0:core_3_mailbox_in_writedata -> core_3:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_4_mailbox_in_readdata;    // core_4:mailbox_in_readdata -> mm_interconnect_0:core_4_mailbox_in_readdata
	wire         mm_interconnect_0_core_4_mailbox_in_waitrequest; // core_4:mailbox_in_waitrequest -> mm_interconnect_0:core_4_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_4_mailbox_in_address;     // mm_interconnect_0:core_4_mailbox_in_address -> core_4:mailbox_in_address
	wire         mm_interconnect_0_core_4_mailbox_in_read;        // mm_interconnect_0:core_4_mailbox_in_read -> core_4:mailbox_in_read
	wire         mm_interconnect_0_core_4_mailbox_in_write;       // mm_interconnect_0:core_4_mailbox_in_write -> core_4:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_4_mailbox_in_writedata;   // mm_interconnect_0:core_4_mailbox_in_writedata -> core_4:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_5_mailbox_in_readdata;    // core_5:mailbox_in_readdata -> mm_interconnect_0:core_5_mailbox_in_readdata
	wire         mm_interconnect_0_core_5_mailbox_in_waitrequest; // core_5:mailbox_in_waitrequest -> mm_interconnect_0:core_5_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_5_mailbox_in_address;     // mm_interconnect_0:core_5_mailbox_in_address -> core_5:mailbox_in_address
	wire         mm_interconnect_0_core_5_mailbox_in_read;        // mm_interconnect_0:core_5_mailbox_in_read -> core_5:mailbox_in_read
	wire         mm_interconnect_0_core_5_mailbox_in_write;       // mm_interconnect_0:core_5_mailbox_in_write -> core_5:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_5_mailbox_in_writedata;   // mm_interconnect_0:core_5_mailbox_in_writedata -> core_5:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_6_mailbox_in_readdata;    // core_6:mailbox_in_readdata -> mm_interconnect_0:core_6_mailbox_in_readdata
	wire         mm_interconnect_0_core_6_mailbox_in_waitrequest; // core_6:mailbox_in_waitrequest -> mm_interconnect_0:core_6_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_6_mailbox_in_address;     // mm_interconnect_0:core_6_mailbox_in_address -> core_6:mailbox_in_address
	wire         mm_interconnect_0_core_6_mailbox_in_read;        // mm_interconnect_0:core_6_mailbox_in_read -> core_6:mailbox_in_read
	wire         mm_interconnect_0_core_6_mailbox_in_write;       // mm_interconnect_0:core_6_mailbox_in_write -> core_6:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_6_mailbox_in_writedata;   // mm_interconnect_0:core_6_mailbox_in_writedata -> core_6:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_7_mailbox_in_readdata;    // core_7:mailbox_in_readdata -> mm_interconnect_0:core_7_mailbox_in_readdata
	wire         mm_interconnect_0_core_7_mailbox_in_waitrequest; // core_7:mailbox_in_waitrequest -> mm_interconnect_0:core_7_mailbox_in_waitrequest
	wire   [1:0] mm_interconnect_0_core_7_mailbox_in_address;     // mm_interconnect_0:core_7_mailbox_in_address -> core_7:mailbox_in_address
	wire         mm_interconnect_0_core_7_mailbox_in_read;        // mm_interconnect_0:core_7_mailbox_in_read -> core_7:mailbox_in_read
	wire         mm_interconnect_0_core_7_mailbox_in_write;       // mm_interconnect_0:core_7_mailbox_in_write -> core_7:mailbox_in_write
	wire  [31:0] mm_interconnect_0_core_7_mailbox_in_writedata;   // mm_interconnect_0:core_7_mailbox_in_writedata -> core_7:mailbox_in_writedata
	wire  [31:0] mm_interconnect_0_core_1_mailbox_out_readdata;   // core_1:mailbox_out_readdata -> mm_interconnect_0:core_1_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_1_mailbox_out_address;    // mm_interconnect_0:core_1_mailbox_out_address -> core_1:mailbox_out_address
	wire         mm_interconnect_0_core_1_mailbox_out_read;       // mm_interconnect_0:core_1_mailbox_out_read -> core_1:mailbox_out_read
	wire         mm_interconnect_0_core_1_mailbox_out_write;      // mm_interconnect_0:core_1_mailbox_out_write -> core_1:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_1_mailbox_out_writedata;  // mm_interconnect_0:core_1_mailbox_out_writedata -> core_1:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_2_mailbox_out_readdata;   // core_2:mailbox_out_readdata -> mm_interconnect_0:core_2_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_2_mailbox_out_address;    // mm_interconnect_0:core_2_mailbox_out_address -> core_2:mailbox_out_address
	wire         mm_interconnect_0_core_2_mailbox_out_read;       // mm_interconnect_0:core_2_mailbox_out_read -> core_2:mailbox_out_read
	wire         mm_interconnect_0_core_2_mailbox_out_write;      // mm_interconnect_0:core_2_mailbox_out_write -> core_2:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_2_mailbox_out_writedata;  // mm_interconnect_0:core_2_mailbox_out_writedata -> core_2:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_3_mailbox_out_readdata;   // core_3:mailbox_out_readdata -> mm_interconnect_0:core_3_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_3_mailbox_out_address;    // mm_interconnect_0:core_3_mailbox_out_address -> core_3:mailbox_out_address
	wire         mm_interconnect_0_core_3_mailbox_out_read;       // mm_interconnect_0:core_3_mailbox_out_read -> core_3:mailbox_out_read
	wire         mm_interconnect_0_core_3_mailbox_out_write;      // mm_interconnect_0:core_3_mailbox_out_write -> core_3:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_3_mailbox_out_writedata;  // mm_interconnect_0:core_3_mailbox_out_writedata -> core_3:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_4_mailbox_out_readdata;   // core_4:mailbox_out_readdata -> mm_interconnect_0:core_4_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_4_mailbox_out_address;    // mm_interconnect_0:core_4_mailbox_out_address -> core_4:mailbox_out_address
	wire         mm_interconnect_0_core_4_mailbox_out_read;       // mm_interconnect_0:core_4_mailbox_out_read -> core_4:mailbox_out_read
	wire         mm_interconnect_0_core_4_mailbox_out_write;      // mm_interconnect_0:core_4_mailbox_out_write -> core_4:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_4_mailbox_out_writedata;  // mm_interconnect_0:core_4_mailbox_out_writedata -> core_4:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_5_mailbox_out_readdata;   // core_5:mailbox_out_readdata -> mm_interconnect_0:core_5_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_5_mailbox_out_address;    // mm_interconnect_0:core_5_mailbox_out_address -> core_5:mailbox_out_address
	wire         mm_interconnect_0_core_5_mailbox_out_read;       // mm_interconnect_0:core_5_mailbox_out_read -> core_5:mailbox_out_read
	wire         mm_interconnect_0_core_5_mailbox_out_write;      // mm_interconnect_0:core_5_mailbox_out_write -> core_5:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_5_mailbox_out_writedata;  // mm_interconnect_0:core_5_mailbox_out_writedata -> core_5:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_6_mailbox_out_readdata;   // core_6:mailbox_out_readdata -> mm_interconnect_0:core_6_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_6_mailbox_out_address;    // mm_interconnect_0:core_6_mailbox_out_address -> core_6:mailbox_out_address
	wire         mm_interconnect_0_core_6_mailbox_out_read;       // mm_interconnect_0:core_6_mailbox_out_read -> core_6:mailbox_out_read
	wire         mm_interconnect_0_core_6_mailbox_out_write;      // mm_interconnect_0:core_6_mailbox_out_write -> core_6:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_6_mailbox_out_writedata;  // mm_interconnect_0:core_6_mailbox_out_writedata -> core_6:mailbox_out_writedata
	wire  [31:0] mm_interconnect_0_core_7_mailbox_out_readdata;   // core_7:mailbox_out_readdata -> mm_interconnect_0:core_7_mailbox_out_readdata
	wire   [1:0] mm_interconnect_0_core_7_mailbox_out_address;    // mm_interconnect_0:core_7_mailbox_out_address -> core_7:mailbox_out_address
	wire         mm_interconnect_0_core_7_mailbox_out_read;       // mm_interconnect_0:core_7_mailbox_out_read -> core_7:mailbox_out_read
	wire         mm_interconnect_0_core_7_mailbox_out_write;      // mm_interconnect_0:core_7_mailbox_out_write -> core_7:mailbox_out_write
	wire  [31:0] mm_interconnect_0_core_7_mailbox_out_writedata;  // mm_interconnect_0:core_7_mailbox_out_writedata -> core_7:mailbox_out_writedata
	wire         mm_interconnect_0_timer_s1_chipselect;           // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;             // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;              // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;            // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_shared_memory_s1_chipselect;   // mm_interconnect_0:shared_memory_s1_chipselect -> shared_memory:chipselect
	wire  [31:0] mm_interconnect_0_shared_memory_s1_readdata;     // shared_memory:readdata -> mm_interconnect_0:shared_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_shared_memory_s1_address;      // mm_interconnect_0:shared_memory_s1_address -> shared_memory:address
	wire   [3:0] mm_interconnect_0_shared_memory_s1_byteenable;   // mm_interconnect_0:shared_memory_s1_byteenable -> shared_memory:byteenable
	wire         mm_interconnect_0_shared_memory_s1_write;        // mm_interconnect_0:shared_memory_s1_write -> shared_memory:write
	wire  [31:0] mm_interconnect_0_shared_memory_s1_writedata;    // mm_interconnect_0:shared_memory_s1_writedata -> shared_memory:writedata
	wire         mm_interconnect_0_shared_memory_s1_clken;        // mm_interconnect_0:shared_memory_s1_clken -> shared_memory:clken
	wire         rst_controller_reset_out_reset;                  // rst_controller:reset_out -> [mm_interconnect_0:core_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, shared_memory:reset, sysid:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;              // rst_controller:reset_req -> [rst_translator:reset_req_in, shared_memory:reset_req]

	multicore_system_core_0 core_0 (
		.clk_clk                   (clk_clk),                          //         clk.clk
		.data_master_waitrequest   (core_0_data_master_waitrequest),   // data_master.waitrequest
		.data_master_readdata      (core_0_data_master_readdata),      //            .readdata
		.data_master_readdatavalid (core_0_data_master_readdatavalid), //            .readdatavalid
		.data_master_burstcount    (core_0_data_master_burstcount),    //            .burstcount
		.data_master_writedata     (core_0_data_master_writedata),     //            .writedata
		.data_master_address       (core_0_data_master_address),       //            .address
		.data_master_write         (core_0_data_master_write),         //            .write
		.data_master_read          (core_0_data_master_read),          //            .read
		.data_master_byteenable    (core_0_data_master_byteenable),    //            .byteenable
		.data_master_debugaccess   (core_0_data_master_debugaccess),   //            .debugaccess
		.mailbox_in_address        (),                                 //  mailbox_in.address
		.mailbox_in_writedata      (),                                 //            .writedata
		.mailbox_in_write          (),                                 //            .write
		.mailbox_in_read           (),                                 //            .read
		.mailbox_in_readdata       (),                                 //            .readdata
		.mailbox_in_waitrequest    (),                                 //            .waitrequest
		.mailbox_out_address       (),                                 // mailbox_out.address
		.mailbox_out_read          (),                                 //            .read
		.mailbox_out_writedata     (),                                 //            .writedata
		.mailbox_out_write         (),                                 //            .write
		.mailbox_out_readdata      (),                                 //            .readdata
		.reset_reset_n             (reset_reset_n)                     //       reset.reset_n
	);

	multicore_system_core_1 core_1 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_1_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_1_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_1_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_1_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_1_data_master_writedata),                    //            .writedata
		.data_master_address       (core_1_data_master_address),                      //            .address
		.data_master_write         (core_1_data_master_write),                        //            .write
		.data_master_read          (core_1_data_master_read),                         //            .read
		.data_master_byteenable    (core_1_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_1_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_1_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_1_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_1_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_1_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_1_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_1_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_1_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_1_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_1_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_1_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_1_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_2 core_2 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_2_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_2_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_2_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_2_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_2_data_master_writedata),                    //            .writedata
		.data_master_address       (core_2_data_master_address),                      //            .address
		.data_master_write         (core_2_data_master_write),                        //            .write
		.data_master_read          (core_2_data_master_read),                         //            .read
		.data_master_byteenable    (core_2_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_2_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_2_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_2_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_2_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_2_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_2_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_2_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_2_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_2_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_2_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_2_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_2_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_3 core_3 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_3_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_3_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_3_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_3_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_3_data_master_writedata),                    //            .writedata
		.data_master_address       (core_3_data_master_address),                      //            .address
		.data_master_write         (core_3_data_master_write),                        //            .write
		.data_master_read          (core_3_data_master_read),                         //            .read
		.data_master_byteenable    (core_3_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_3_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_3_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_3_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_3_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_3_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_3_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_3_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_3_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_3_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_3_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_3_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_3_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_4 core_4 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_4_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_4_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_4_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_4_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_4_data_master_writedata),                    //            .writedata
		.data_master_address       (core_4_data_master_address),                      //            .address
		.data_master_write         (core_4_data_master_write),                        //            .write
		.data_master_read          (core_4_data_master_read),                         //            .read
		.data_master_byteenable    (core_4_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_4_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_4_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_4_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_4_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_4_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_4_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_4_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_4_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_4_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_4_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_4_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_4_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_5 core_5 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_5_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_5_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_5_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_5_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_5_data_master_writedata),                    //            .writedata
		.data_master_address       (core_5_data_master_address),                      //            .address
		.data_master_write         (core_5_data_master_write),                        //            .write
		.data_master_read          (core_5_data_master_read),                         //            .read
		.data_master_byteenable    (core_5_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_5_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_5_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_5_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_5_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_5_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_5_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_5_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_5_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_5_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_5_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_5_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_5_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_6 core_6 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_6_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_6_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_6_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_6_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_6_data_master_writedata),                    //            .writedata
		.data_master_address       (core_6_data_master_address),                      //            .address
		.data_master_write         (core_6_data_master_write),                        //            .write
		.data_master_read          (core_6_data_master_read),                         //            .read
		.data_master_byteenable    (core_6_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_6_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_6_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_6_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_6_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_6_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_6_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_6_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_6_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_6_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_6_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_6_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_6_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_core_7 core_7 (
		.clk_clk                   (clk_clk),                                         //         clk.clk
		.data_master_waitrequest   (core_7_data_master_waitrequest),                  // data_master.waitrequest
		.data_master_readdata      (core_7_data_master_readdata),                     //            .readdata
		.data_master_readdatavalid (core_7_data_master_readdatavalid),                //            .readdatavalid
		.data_master_burstcount    (core_7_data_master_burstcount),                   //            .burstcount
		.data_master_writedata     (core_7_data_master_writedata),                    //            .writedata
		.data_master_address       (core_7_data_master_address),                      //            .address
		.data_master_write         (core_7_data_master_write),                        //            .write
		.data_master_read          (core_7_data_master_read),                         //            .read
		.data_master_byteenable    (core_7_data_master_byteenable),                   //            .byteenable
		.data_master_debugaccess   (core_7_data_master_debugaccess),                  //            .debugaccess
		.mailbox_in_address        (mm_interconnect_0_core_7_mailbox_in_address),     //  mailbox_in.address
		.mailbox_in_writedata      (mm_interconnect_0_core_7_mailbox_in_writedata),   //            .writedata
		.mailbox_in_write          (mm_interconnect_0_core_7_mailbox_in_write),       //            .write
		.mailbox_in_read           (mm_interconnect_0_core_7_mailbox_in_read),        //            .read
		.mailbox_in_readdata       (mm_interconnect_0_core_7_mailbox_in_readdata),    //            .readdata
		.mailbox_in_waitrequest    (mm_interconnect_0_core_7_mailbox_in_waitrequest), //            .waitrequest
		.mailbox_out_address       (mm_interconnect_0_core_7_mailbox_out_address),    // mailbox_out.address
		.mailbox_out_read          (mm_interconnect_0_core_7_mailbox_out_read),       //            .read
		.mailbox_out_writedata     (mm_interconnect_0_core_7_mailbox_out_writedata),  //            .writedata
		.mailbox_out_write         (mm_interconnect_0_core_7_mailbox_out_write),      //            .write
		.mailbox_out_readdata      (mm_interconnect_0_core_7_mailbox_out_readdata),   //            .readdata
		.reset_reset_n             (reset_reset_n)                                    //       reset.reset_n
	);

	multicore_system_shared_memory shared_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_shared_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_shared_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_shared_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_shared_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_shared_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_shared_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_shared_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	multicore_system_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	multicore_system_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        ()                                       //   irq.irq
	);

	multicore_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (clk_clk),                                         //                            clk_clk.clk
		.core_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                  // core_0_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                  //  sysid_reset_reset_bridge_in_reset.reset
		.core_0_data_master_address               (core_0_data_master_address),                      //                 core_0_data_master.address
		.core_0_data_master_waitrequest           (core_0_data_master_waitrequest),                  //                                   .waitrequest
		.core_0_data_master_burstcount            (core_0_data_master_burstcount),                   //                                   .burstcount
		.core_0_data_master_byteenable            (core_0_data_master_byteenable),                   //                                   .byteenable
		.core_0_data_master_read                  (core_0_data_master_read),                         //                                   .read
		.core_0_data_master_readdata              (core_0_data_master_readdata),                     //                                   .readdata
		.core_0_data_master_readdatavalid         (core_0_data_master_readdatavalid),                //                                   .readdatavalid
		.core_0_data_master_write                 (core_0_data_master_write),                        //                                   .write
		.core_0_data_master_writedata             (core_0_data_master_writedata),                    //                                   .writedata
		.core_0_data_master_debugaccess           (core_0_data_master_debugaccess),                  //                                   .debugaccess
		.core_1_data_master_address               (core_1_data_master_address),                      //                 core_1_data_master.address
		.core_1_data_master_waitrequest           (core_1_data_master_waitrequest),                  //                                   .waitrequest
		.core_1_data_master_burstcount            (core_1_data_master_burstcount),                   //                                   .burstcount
		.core_1_data_master_byteenable            (core_1_data_master_byteenable),                   //                                   .byteenable
		.core_1_data_master_read                  (core_1_data_master_read),                         //                                   .read
		.core_1_data_master_readdata              (core_1_data_master_readdata),                     //                                   .readdata
		.core_1_data_master_readdatavalid         (core_1_data_master_readdatavalid),                //                                   .readdatavalid
		.core_1_data_master_write                 (core_1_data_master_write),                        //                                   .write
		.core_1_data_master_writedata             (core_1_data_master_writedata),                    //                                   .writedata
		.core_1_data_master_debugaccess           (core_1_data_master_debugaccess),                  //                                   .debugaccess
		.core_2_data_master_address               (core_2_data_master_address),                      //                 core_2_data_master.address
		.core_2_data_master_waitrequest           (core_2_data_master_waitrequest),                  //                                   .waitrequest
		.core_2_data_master_burstcount            (core_2_data_master_burstcount),                   //                                   .burstcount
		.core_2_data_master_byteenable            (core_2_data_master_byteenable),                   //                                   .byteenable
		.core_2_data_master_read                  (core_2_data_master_read),                         //                                   .read
		.core_2_data_master_readdata              (core_2_data_master_readdata),                     //                                   .readdata
		.core_2_data_master_readdatavalid         (core_2_data_master_readdatavalid),                //                                   .readdatavalid
		.core_2_data_master_write                 (core_2_data_master_write),                        //                                   .write
		.core_2_data_master_writedata             (core_2_data_master_writedata),                    //                                   .writedata
		.core_2_data_master_debugaccess           (core_2_data_master_debugaccess),                  //                                   .debugaccess
		.core_3_data_master_address               (core_3_data_master_address),                      //                 core_3_data_master.address
		.core_3_data_master_waitrequest           (core_3_data_master_waitrequest),                  //                                   .waitrequest
		.core_3_data_master_burstcount            (core_3_data_master_burstcount),                   //                                   .burstcount
		.core_3_data_master_byteenable            (core_3_data_master_byteenable),                   //                                   .byteenable
		.core_3_data_master_read                  (core_3_data_master_read),                         //                                   .read
		.core_3_data_master_readdata              (core_3_data_master_readdata),                     //                                   .readdata
		.core_3_data_master_readdatavalid         (core_3_data_master_readdatavalid),                //                                   .readdatavalid
		.core_3_data_master_write                 (core_3_data_master_write),                        //                                   .write
		.core_3_data_master_writedata             (core_3_data_master_writedata),                    //                                   .writedata
		.core_3_data_master_debugaccess           (core_3_data_master_debugaccess),                  //                                   .debugaccess
		.core_4_data_master_address               (core_4_data_master_address),                      //                 core_4_data_master.address
		.core_4_data_master_waitrequest           (core_4_data_master_waitrequest),                  //                                   .waitrequest
		.core_4_data_master_burstcount            (core_4_data_master_burstcount),                   //                                   .burstcount
		.core_4_data_master_byteenable            (core_4_data_master_byteenable),                   //                                   .byteenable
		.core_4_data_master_read                  (core_4_data_master_read),                         //                                   .read
		.core_4_data_master_readdata              (core_4_data_master_readdata),                     //                                   .readdata
		.core_4_data_master_readdatavalid         (core_4_data_master_readdatavalid),                //                                   .readdatavalid
		.core_4_data_master_write                 (core_4_data_master_write),                        //                                   .write
		.core_4_data_master_writedata             (core_4_data_master_writedata),                    //                                   .writedata
		.core_4_data_master_debugaccess           (core_4_data_master_debugaccess),                  //                                   .debugaccess
		.core_5_data_master_address               (core_5_data_master_address),                      //                 core_5_data_master.address
		.core_5_data_master_waitrequest           (core_5_data_master_waitrequest),                  //                                   .waitrequest
		.core_5_data_master_burstcount            (core_5_data_master_burstcount),                   //                                   .burstcount
		.core_5_data_master_byteenable            (core_5_data_master_byteenable),                   //                                   .byteenable
		.core_5_data_master_read                  (core_5_data_master_read),                         //                                   .read
		.core_5_data_master_readdata              (core_5_data_master_readdata),                     //                                   .readdata
		.core_5_data_master_readdatavalid         (core_5_data_master_readdatavalid),                //                                   .readdatavalid
		.core_5_data_master_write                 (core_5_data_master_write),                        //                                   .write
		.core_5_data_master_writedata             (core_5_data_master_writedata),                    //                                   .writedata
		.core_5_data_master_debugaccess           (core_5_data_master_debugaccess),                  //                                   .debugaccess
		.core_6_data_master_address               (core_6_data_master_address),                      //                 core_6_data_master.address
		.core_6_data_master_waitrequest           (core_6_data_master_waitrequest),                  //                                   .waitrequest
		.core_6_data_master_burstcount            (core_6_data_master_burstcount),                   //                                   .burstcount
		.core_6_data_master_byteenable            (core_6_data_master_byteenable),                   //                                   .byteenable
		.core_6_data_master_read                  (core_6_data_master_read),                         //                                   .read
		.core_6_data_master_readdata              (core_6_data_master_readdata),                     //                                   .readdata
		.core_6_data_master_readdatavalid         (core_6_data_master_readdatavalid),                //                                   .readdatavalid
		.core_6_data_master_write                 (core_6_data_master_write),                        //                                   .write
		.core_6_data_master_writedata             (core_6_data_master_writedata),                    //                                   .writedata
		.core_6_data_master_debugaccess           (core_6_data_master_debugaccess),                  //                                   .debugaccess
		.core_7_data_master_address               (core_7_data_master_address),                      //                 core_7_data_master.address
		.core_7_data_master_waitrequest           (core_7_data_master_waitrequest),                  //                                   .waitrequest
		.core_7_data_master_burstcount            (core_7_data_master_burstcount),                   //                                   .burstcount
		.core_7_data_master_byteenable            (core_7_data_master_byteenable),                   //                                   .byteenable
		.core_7_data_master_read                  (core_7_data_master_read),                         //                                   .read
		.core_7_data_master_readdata              (core_7_data_master_readdata),                     //                                   .readdata
		.core_7_data_master_readdatavalid         (core_7_data_master_readdatavalid),                //                                   .readdatavalid
		.core_7_data_master_write                 (core_7_data_master_write),                        //                                   .write
		.core_7_data_master_writedata             (core_7_data_master_writedata),                    //                                   .writedata
		.core_7_data_master_debugaccess           (core_7_data_master_debugaccess),                  //                                   .debugaccess
		.core_1_mailbox_in_address                (mm_interconnect_0_core_1_mailbox_in_address),     //                  core_1_mailbox_in.address
		.core_1_mailbox_in_write                  (mm_interconnect_0_core_1_mailbox_in_write),       //                                   .write
		.core_1_mailbox_in_read                   (mm_interconnect_0_core_1_mailbox_in_read),        //                                   .read
		.core_1_mailbox_in_readdata               (mm_interconnect_0_core_1_mailbox_in_readdata),    //                                   .readdata
		.core_1_mailbox_in_writedata              (mm_interconnect_0_core_1_mailbox_in_writedata),   //                                   .writedata
		.core_1_mailbox_in_waitrequest            (mm_interconnect_0_core_1_mailbox_in_waitrequest), //                                   .waitrequest
		.core_1_mailbox_out_address               (mm_interconnect_0_core_1_mailbox_out_address),    //                 core_1_mailbox_out.address
		.core_1_mailbox_out_write                 (mm_interconnect_0_core_1_mailbox_out_write),      //                                   .write
		.core_1_mailbox_out_read                  (mm_interconnect_0_core_1_mailbox_out_read),       //                                   .read
		.core_1_mailbox_out_readdata              (mm_interconnect_0_core_1_mailbox_out_readdata),   //                                   .readdata
		.core_1_mailbox_out_writedata             (mm_interconnect_0_core_1_mailbox_out_writedata),  //                                   .writedata
		.core_2_mailbox_in_address                (mm_interconnect_0_core_2_mailbox_in_address),     //                  core_2_mailbox_in.address
		.core_2_mailbox_in_write                  (mm_interconnect_0_core_2_mailbox_in_write),       //                                   .write
		.core_2_mailbox_in_read                   (mm_interconnect_0_core_2_mailbox_in_read),        //                                   .read
		.core_2_mailbox_in_readdata               (mm_interconnect_0_core_2_mailbox_in_readdata),    //                                   .readdata
		.core_2_mailbox_in_writedata              (mm_interconnect_0_core_2_mailbox_in_writedata),   //                                   .writedata
		.core_2_mailbox_in_waitrequest            (mm_interconnect_0_core_2_mailbox_in_waitrequest), //                                   .waitrequest
		.core_2_mailbox_out_address               (mm_interconnect_0_core_2_mailbox_out_address),    //                 core_2_mailbox_out.address
		.core_2_mailbox_out_write                 (mm_interconnect_0_core_2_mailbox_out_write),      //                                   .write
		.core_2_mailbox_out_read                  (mm_interconnect_0_core_2_mailbox_out_read),       //                                   .read
		.core_2_mailbox_out_readdata              (mm_interconnect_0_core_2_mailbox_out_readdata),   //                                   .readdata
		.core_2_mailbox_out_writedata             (mm_interconnect_0_core_2_mailbox_out_writedata),  //                                   .writedata
		.core_3_mailbox_in_address                (mm_interconnect_0_core_3_mailbox_in_address),     //                  core_3_mailbox_in.address
		.core_3_mailbox_in_write                  (mm_interconnect_0_core_3_mailbox_in_write),       //                                   .write
		.core_3_mailbox_in_read                   (mm_interconnect_0_core_3_mailbox_in_read),        //                                   .read
		.core_3_mailbox_in_readdata               (mm_interconnect_0_core_3_mailbox_in_readdata),    //                                   .readdata
		.core_3_mailbox_in_writedata              (mm_interconnect_0_core_3_mailbox_in_writedata),   //                                   .writedata
		.core_3_mailbox_in_waitrequest            (mm_interconnect_0_core_3_mailbox_in_waitrequest), //                                   .waitrequest
		.core_3_mailbox_out_address               (mm_interconnect_0_core_3_mailbox_out_address),    //                 core_3_mailbox_out.address
		.core_3_mailbox_out_write                 (mm_interconnect_0_core_3_mailbox_out_write),      //                                   .write
		.core_3_mailbox_out_read                  (mm_interconnect_0_core_3_mailbox_out_read),       //                                   .read
		.core_3_mailbox_out_readdata              (mm_interconnect_0_core_3_mailbox_out_readdata),   //                                   .readdata
		.core_3_mailbox_out_writedata             (mm_interconnect_0_core_3_mailbox_out_writedata),  //                                   .writedata
		.core_4_mailbox_in_address                (mm_interconnect_0_core_4_mailbox_in_address),     //                  core_4_mailbox_in.address
		.core_4_mailbox_in_write                  (mm_interconnect_0_core_4_mailbox_in_write),       //                                   .write
		.core_4_mailbox_in_read                   (mm_interconnect_0_core_4_mailbox_in_read),        //                                   .read
		.core_4_mailbox_in_readdata               (mm_interconnect_0_core_4_mailbox_in_readdata),    //                                   .readdata
		.core_4_mailbox_in_writedata              (mm_interconnect_0_core_4_mailbox_in_writedata),   //                                   .writedata
		.core_4_mailbox_in_waitrequest            (mm_interconnect_0_core_4_mailbox_in_waitrequest), //                                   .waitrequest
		.core_4_mailbox_out_address               (mm_interconnect_0_core_4_mailbox_out_address),    //                 core_4_mailbox_out.address
		.core_4_mailbox_out_write                 (mm_interconnect_0_core_4_mailbox_out_write),      //                                   .write
		.core_4_mailbox_out_read                  (mm_interconnect_0_core_4_mailbox_out_read),       //                                   .read
		.core_4_mailbox_out_readdata              (mm_interconnect_0_core_4_mailbox_out_readdata),   //                                   .readdata
		.core_4_mailbox_out_writedata             (mm_interconnect_0_core_4_mailbox_out_writedata),  //                                   .writedata
		.core_5_mailbox_in_address                (mm_interconnect_0_core_5_mailbox_in_address),     //                  core_5_mailbox_in.address
		.core_5_mailbox_in_write                  (mm_interconnect_0_core_5_mailbox_in_write),       //                                   .write
		.core_5_mailbox_in_read                   (mm_interconnect_0_core_5_mailbox_in_read),        //                                   .read
		.core_5_mailbox_in_readdata               (mm_interconnect_0_core_5_mailbox_in_readdata),    //                                   .readdata
		.core_5_mailbox_in_writedata              (mm_interconnect_0_core_5_mailbox_in_writedata),   //                                   .writedata
		.core_5_mailbox_in_waitrequest            (mm_interconnect_0_core_5_mailbox_in_waitrequest), //                                   .waitrequest
		.core_5_mailbox_out_address               (mm_interconnect_0_core_5_mailbox_out_address),    //                 core_5_mailbox_out.address
		.core_5_mailbox_out_write                 (mm_interconnect_0_core_5_mailbox_out_write),      //                                   .write
		.core_5_mailbox_out_read                  (mm_interconnect_0_core_5_mailbox_out_read),       //                                   .read
		.core_5_mailbox_out_readdata              (mm_interconnect_0_core_5_mailbox_out_readdata),   //                                   .readdata
		.core_5_mailbox_out_writedata             (mm_interconnect_0_core_5_mailbox_out_writedata),  //                                   .writedata
		.core_6_mailbox_in_address                (mm_interconnect_0_core_6_mailbox_in_address),     //                  core_6_mailbox_in.address
		.core_6_mailbox_in_write                  (mm_interconnect_0_core_6_mailbox_in_write),       //                                   .write
		.core_6_mailbox_in_read                   (mm_interconnect_0_core_6_mailbox_in_read),        //                                   .read
		.core_6_mailbox_in_readdata               (mm_interconnect_0_core_6_mailbox_in_readdata),    //                                   .readdata
		.core_6_mailbox_in_writedata              (mm_interconnect_0_core_6_mailbox_in_writedata),   //                                   .writedata
		.core_6_mailbox_in_waitrequest            (mm_interconnect_0_core_6_mailbox_in_waitrequest), //                                   .waitrequest
		.core_6_mailbox_out_address               (mm_interconnect_0_core_6_mailbox_out_address),    //                 core_6_mailbox_out.address
		.core_6_mailbox_out_write                 (mm_interconnect_0_core_6_mailbox_out_write),      //                                   .write
		.core_6_mailbox_out_read                  (mm_interconnect_0_core_6_mailbox_out_read),       //                                   .read
		.core_6_mailbox_out_readdata              (mm_interconnect_0_core_6_mailbox_out_readdata),   //                                   .readdata
		.core_6_mailbox_out_writedata             (mm_interconnect_0_core_6_mailbox_out_writedata),  //                                   .writedata
		.core_7_mailbox_in_address                (mm_interconnect_0_core_7_mailbox_in_address),     //                  core_7_mailbox_in.address
		.core_7_mailbox_in_write                  (mm_interconnect_0_core_7_mailbox_in_write),       //                                   .write
		.core_7_mailbox_in_read                   (mm_interconnect_0_core_7_mailbox_in_read),        //                                   .read
		.core_7_mailbox_in_readdata               (mm_interconnect_0_core_7_mailbox_in_readdata),    //                                   .readdata
		.core_7_mailbox_in_writedata              (mm_interconnect_0_core_7_mailbox_in_writedata),   //                                   .writedata
		.core_7_mailbox_in_waitrequest            (mm_interconnect_0_core_7_mailbox_in_waitrequest), //                                   .waitrequest
		.core_7_mailbox_out_address               (mm_interconnect_0_core_7_mailbox_out_address),    //                 core_7_mailbox_out.address
		.core_7_mailbox_out_write                 (mm_interconnect_0_core_7_mailbox_out_write),      //                                   .write
		.core_7_mailbox_out_read                  (mm_interconnect_0_core_7_mailbox_out_read),       //                                   .read
		.core_7_mailbox_out_readdata              (mm_interconnect_0_core_7_mailbox_out_readdata),   //                                   .readdata
		.core_7_mailbox_out_writedata             (mm_interconnect_0_core_7_mailbox_out_writedata),  //                                   .writedata
		.shared_memory_s1_address                 (mm_interconnect_0_shared_memory_s1_address),      //                   shared_memory_s1.address
		.shared_memory_s1_write                   (mm_interconnect_0_shared_memory_s1_write),        //                                   .write
		.shared_memory_s1_readdata                (mm_interconnect_0_shared_memory_s1_readdata),     //                                   .readdata
		.shared_memory_s1_writedata               (mm_interconnect_0_shared_memory_s1_writedata),    //                                   .writedata
		.shared_memory_s1_byteenable              (mm_interconnect_0_shared_memory_s1_byteenable),   //                                   .byteenable
		.shared_memory_s1_chipselect              (mm_interconnect_0_shared_memory_s1_chipselect),   //                                   .chipselect
		.shared_memory_s1_clken                   (mm_interconnect_0_shared_memory_s1_clken),        //                                   .clken
		.sysid_control_slave_address              (mm_interconnect_0_sysid_control_slave_address),   //                sysid_control_slave.address
		.sysid_control_slave_readdata             (mm_interconnect_0_sysid_control_slave_readdata),  //                                   .readdata
		.timer_s1_address                         (mm_interconnect_0_timer_s1_address),              //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_0_timer_s1_write),                //                                   .write
		.timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),             //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),            //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect)            //                                   .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
