// multicore_system_core_3.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module multicore_system_core_3 (
		input  wire        clk_clk,                   //         clk.clk
		input  wire        data_master_waitrequest,   // data_master.waitrequest
		input  wire [31:0] data_master_readdata,      //            .readdata
		input  wire        data_master_readdatavalid, //            .readdatavalid
		output wire [0:0]  data_master_burstcount,    //            .burstcount
		output wire [31:0] data_master_writedata,     //            .writedata
		output wire [19:0] data_master_address,       //            .address
		output wire        data_master_write,         //            .write
		output wire        data_master_read,          //            .read
		output wire [3:0]  data_master_byteenable,    //            .byteenable
		output wire        data_master_debugaccess,   //            .debugaccess
		input  wire [1:0]  mailbox_in_address,        //  mailbox_in.address
		input  wire [31:0] mailbox_in_writedata,      //            .writedata
		input  wire        mailbox_in_write,          //            .write
		input  wire        mailbox_in_read,           //            .read
		output wire [31:0] mailbox_in_readdata,       //            .readdata
		output wire        mailbox_in_waitrequest,    //            .waitrequest
		input  wire [1:0]  mailbox_out_address,       // mailbox_out.address
		input  wire        mailbox_out_read,          //            .read
		input  wire [31:0] mailbox_out_writedata,     //            .writedata
		input  wire        mailbox_out_write,         //            .write
		output wire [31:0] mailbox_out_readdata,      //            .readdata
		input  wire        reset_reset_n              //       reset.reset_n
	);

	wire  [31:0] nios2_custom_instruction_master_multi_dataa;                              // nios2:A_ci_multi_dataa -> nios2_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_custom_instruction_master_multi_writerc;                            // nios2:A_ci_multi_writerc -> nios2_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_result;                             // nios2_custom_instruction_master_translator:ci_slave_multi_result -> nios2:A_ci_multi_result
	wire         nios2_custom_instruction_master_clk;                                      // nios2:A_ci_multi_clock -> nios2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_custom_instruction_master_multi_datab;                              // nios2:A_ci_multi_datab -> nios2_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_custom_instruction_master_start;                                    // nios2:A_ci_multi_start -> nios2_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_custom_instruction_master_multi_b;                                  // nios2:A_ci_multi_b -> nios2_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_custom_instruction_master_multi_c;                                  // nios2:A_ci_multi_c -> nios2_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_custom_instruction_master_reset_req;                                // nios2:A_ci_multi_reset_req -> nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_custom_instruction_master_done;                                     // nios2_custom_instruction_master_translator:ci_slave_multi_done -> nios2:A_ci_multi_done
	wire   [4:0] nios2_custom_instruction_master_multi_a;                                  // nios2:A_ci_multi_a -> nios2_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_custom_instruction_master_clk_en;                                   // nios2:A_ci_multi_clk_en -> nios2_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_custom_instruction_master_reset;                                    // nios2:A_ci_multi_reset -> nios2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_custom_instruction_master_multi_readrb;                             // nios2:A_ci_multi_readrb -> nios2_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_custom_instruction_master_multi_readra;                             // nios2:A_ci_multi_readra -> nios2_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_custom_instruction_master_multi_n;                                  // nios2:A_ci_multi_n -> nios2_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_custom_instruction_master_translator:multi_ci_master_readra -> nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_a;             // nios2_custom_instruction_master_translator:multi_ci_master_a -> nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_b;             // nios2_custom_instruction_master_translator:multi_ci_master_b -> nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_custom_instruction_master_translator:multi_ci_master_clk -> nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_c;             // nios2_custom_instruction_master_translator:multi_ci_master_c -> nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_custom_instruction_master_translator_multi_ci_master_start;         // nios2_custom_instruction_master_translator:multi_ci_master_start -> nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_custom_instruction_master_translator_multi_ci_master_done;          // nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_custom_instruction_master_translator_multi_ci_master_n;             // nios2_custom_instruction_master_translator:multi_ci_master_n -> nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_result;        // nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_custom_instruction_master_translator:multi_ci_master_clken -> nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_custom_instruction_master_translator:multi_ci_master_datab -> nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_custom_instruction_master_translator:multi_ci_master_reset -> nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_result; // custom_instruction:result -> nios2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> custom_instruction:clk
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> custom_instruction:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> custom_instruction:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> custom_instruction:dataa
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_start -> custom_instruction:start
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> custom_instruction:reset
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_done;   // custom_instruction:done -> nios2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [7:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_n;      // nios2_custom_instruction_master_multi_slave_translator0:ci_master_n -> custom_instruction:n
	wire  [31:0] nios2_data_master_readdata;                                               // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                            // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                            // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [20:0] nios2_data_master_address;                                                // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                             // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                   // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_readdatavalid;                                          // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire         nios2_data_master_write;                                                  // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                              // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire   [3:0] nios2_data_master_burstcount;                                             // nios2:d_burstcount -> mm_interconnect_0:nios2_data_master_burstcount
	wire  [31:0] nios2_instruction_master_readdata;                                        // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [20:0] nios2_instruction_master_address;                                         // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                            // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                      // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                        // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                     // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                         // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                            // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                           // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                       // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_readdata;           // avalon_mailbox_in:avmm_rcv_readdata -> mm_interconnect_0:avalon_mailbox_in_avmm_msg_receiver_readdata
	wire   [1:0] mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_address;            // mm_interconnect_0:avalon_mailbox_in_avmm_msg_receiver_address -> avalon_mailbox_in:avmm_rcv_address
	wire         mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_read;               // mm_interconnect_0:avalon_mailbox_in_avmm_msg_receiver_read -> avalon_mailbox_in:avmm_rcv_read
	wire         mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_write;              // mm_interconnect_0:avalon_mailbox_in_avmm_msg_receiver_write -> avalon_mailbox_in:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_writedata;          // mm_interconnect_0:avalon_mailbox_in_avmm_msg_receiver_writedata -> avalon_mailbox_in:avmm_rcv_writedata
	wire  [31:0] mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_readdata;            // avalon_mailbox_out:avmm_snd_readdata -> mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_readdata
	wire         mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_waitrequest;         // avalon_mailbox_out:avmm_snd_waitrequest -> mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_waitrequest
	wire   [1:0] mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_address;             // mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_address -> avalon_mailbox_out:avmm_snd_address
	wire         mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_read;                // mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_read -> avalon_mailbox_out:avmm_snd_read
	wire         mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_write;               // mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_write -> avalon_mailbox_out:avmm_snd_write
	wire  [31:0] mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_writedata;           // mm_interconnect_0:avalon_mailbox_out_avmm_msg_sender_writedata -> avalon_mailbox_out:avmm_snd_writedata
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                         // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                      // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                          // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                             // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                            // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_avalon_data_bridge_s0_readdata;                         // avalon_data_bridge:s0_readdata -> mm_interconnect_0:avalon_data_bridge_s0_readdata
	wire         mm_interconnect_0_avalon_data_bridge_s0_waitrequest;                      // avalon_data_bridge:s0_waitrequest -> mm_interconnect_0:avalon_data_bridge_s0_waitrequest
	wire         mm_interconnect_0_avalon_data_bridge_s0_debugaccess;                      // mm_interconnect_0:avalon_data_bridge_s0_debugaccess -> avalon_data_bridge:s0_debugaccess
	wire  [19:0] mm_interconnect_0_avalon_data_bridge_s0_address;                          // mm_interconnect_0:avalon_data_bridge_s0_address -> avalon_data_bridge:s0_address
	wire         mm_interconnect_0_avalon_data_bridge_s0_read;                             // mm_interconnect_0:avalon_data_bridge_s0_read -> avalon_data_bridge:s0_read
	wire   [3:0] mm_interconnect_0_avalon_data_bridge_s0_byteenable;                       // mm_interconnect_0:avalon_data_bridge_s0_byteenable -> avalon_data_bridge:s0_byteenable
	wire         mm_interconnect_0_avalon_data_bridge_s0_readdatavalid;                    // avalon_data_bridge:s0_readdatavalid -> mm_interconnect_0:avalon_data_bridge_s0_readdatavalid
	wire         mm_interconnect_0_avalon_data_bridge_s0_write;                            // mm_interconnect_0:avalon_data_bridge_s0_write -> avalon_data_bridge:s0_write
	wire  [31:0] mm_interconnect_0_avalon_data_bridge_s0_writedata;                        // mm_interconnect_0:avalon_data_bridge_s0_writedata -> avalon_data_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_avalon_data_bridge_s0_burstcount;                       // mm_interconnect_0:avalon_data_bridge_s0_burstcount -> avalon_data_bridge:s0_burstcount
	wire         mm_interconnect_0_timer_s1_chipselect;                                    // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                      // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                       // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                         // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                     // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_rom_s2_chipselect;                                      // mm_interconnect_0:rom_s2_chipselect -> rom:chipselect2
	wire  [31:0] mm_interconnect_0_rom_s2_readdata;                                        // rom:readdata2 -> mm_interconnect_0:rom_s2_readdata
	wire  [11:0] mm_interconnect_0_rom_s2_address;                                         // mm_interconnect_0:rom_s2_address -> rom:address2
	wire   [3:0] mm_interconnect_0_rom_s2_byteenable;                                      // mm_interconnect_0:rom_s2_byteenable -> rom:byteenable2
	wire         mm_interconnect_0_rom_s2_write;                                           // mm_interconnect_0:rom_s2_write -> rom:write2
	wire  [31:0] mm_interconnect_0_rom_s2_writedata;                                       // mm_interconnect_0:rom_s2_writedata -> rom:writedata2
	wire         mm_interconnect_0_rom_s2_clken;                                           // mm_interconnect_0:rom_s2_clken -> rom:clken2
	wire  [31:0] nios2_tightly_coupled_data_master_0_readdata;                             // mm_interconnect_1:nios2_tightly_coupled_data_master_0_readdata -> nios2:dtcm0_readdata
	wire  [20:0] nios2_tightly_coupled_data_master_0_address;                              // nios2:dtcm0_address -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_address
	wire         nios2_tightly_coupled_data_master_0_read;                                 // nios2:dtcm0_read -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_read
	wire   [3:0] nios2_tightly_coupled_data_master_0_byteenable;                           // nios2:dtcm0_byteenable -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_byteenable
	wire         nios2_tightly_coupled_data_master_0_write;                                // nios2:dtcm0_write -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_write
	wire  [31:0] nios2_tightly_coupled_data_master_0_writedata;                            // nios2:dtcm0_writedata -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_writedata
	wire         nios2_tightly_coupled_data_master_0_clken;                                // nios2:dtcm0_clken -> mm_interconnect_1:nios2_tightly_coupled_data_master_0_clken
	wire         mm_interconnect_1_ram_s1_chipselect;                                      // mm_interconnect_1:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_1_ram_s1_readdata;                                        // ram:readdata -> mm_interconnect_1:ram_s1_readdata
	wire   [9:0] mm_interconnect_1_ram_s1_address;                                         // mm_interconnect_1:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_1_ram_s1_byteenable;                                      // mm_interconnect_1:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_1_ram_s1_write;                                           // mm_interconnect_1:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_1_ram_s1_writedata;                                       // mm_interconnect_1:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_1_ram_s1_clken;                                           // mm_interconnect_1:ram_s1_clken -> ram:clken
	wire  [31:0] nios2_tightly_coupled_instruction_master_0_readdata;                      // mm_interconnect_2:nios2_tightly_coupled_instruction_master_0_readdata -> nios2:itcm0_readdata
	wire  [20:0] nios2_tightly_coupled_instruction_master_0_address;                       // nios2:itcm0_address -> mm_interconnect_2:nios2_tightly_coupled_instruction_master_0_address
	wire         nios2_tightly_coupled_instruction_master_0_read;                          // nios2:itcm0_read -> mm_interconnect_2:nios2_tightly_coupled_instruction_master_0_read
	wire         nios2_tightly_coupled_instruction_master_0_clken;                         // nios2:itcm0_clken -> mm_interconnect_2:nios2_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_2_rom_s1_chipselect;                                      // mm_interconnect_2:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_2_rom_s1_readdata;                                        // rom:readdata -> mm_interconnect_2:rom_s1_readdata
	wire  [11:0] mm_interconnect_2_rom_s1_address;                                         // mm_interconnect_2:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_2_rom_s1_byteenable;                                      // mm_interconnect_2:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_2_rom_s1_write;                                           // mm_interconnect_2:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_2_rom_s1_writedata;                                       // mm_interconnect_2:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_2_rom_s1_clken;                                           // mm_interconnect_2:rom_s1_clken -> rom:clken
	wire         irq_mapper_receiver0_irq;                                                 // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                 // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                                            // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                                           // rst_controller:reset_out -> [avalon_data_bridge:reset, avalon_mailbox_in:rst_n, avalon_mailbox_out:rst_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_reset_reset_bridge_in_reset_reset, mm_interconnect_2:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, ram:reset, rom:reset, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                       // rst_controller:reset_req -> [nios2:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                                          // nios2:debug_reset_request -> rst_controller:reset_in1

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (20),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) avalon_data_bridge (
		.clk              (clk_clk),                                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                        // reset.reset
		.s0_waitrequest   (mm_interconnect_0_avalon_data_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_avalon_data_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_avalon_data_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_avalon_data_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_avalon_data_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_avalon_data_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_avalon_data_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_avalon_data_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_avalon_data_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_avalon_data_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (data_master_waitrequest),                               //    m0.waitrequest
		.m0_readdata      (data_master_readdata),                                  //      .readdata
		.m0_readdatavalid (data_master_readdatavalid),                             //      .readdatavalid
		.m0_burstcount    (data_master_burstcount),                                //      .burstcount
		.m0_writedata     (data_master_writedata),                                 //      .writedata
		.m0_address       (data_master_address),                                   //      .address
		.m0_write         (data_master_write),                                     //      .write
		.m0_read          (data_master_read),                                      //      .read
		.m0_byteenable    (data_master_byteenable),                                //      .byteenable
		.m0_debugaccess   (data_master_debugaccess),                               //      .debugaccess
		.s0_response      (),                                                      // (terminated)
		.m0_response      (2'b00)                                                  // (terminated)
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) avalon_mailbox_in (
		.clk                  (clk_clk),                                                         //               clk.clk
		.rst_n                (~rst_controller_reset_out_reset),                                 //             rst_n.reset_n
		.avmm_snd_address     (mailbox_in_address),                                              //   avmm_msg_sender.address
		.avmm_snd_writedata   (mailbox_in_writedata),                                            //                  .writedata
		.avmm_snd_write       (mailbox_in_write),                                                //                  .write
		.avmm_snd_read        (mailbox_in_read),                                                 //                  .read
		.avmm_snd_readdata    (mailbox_in_readdata),                                             //                  .readdata
		.avmm_snd_waitrequest (mailbox_in_waitrequest),                                          //                  .waitrequest
		.avmm_rcv_address     (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_address),   // avmm_msg_receiver.address
		.avmm_rcv_read        (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_read),      //                  .read
		.avmm_rcv_writedata   (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_writedata), //                  .writedata
		.avmm_rcv_write       (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_write),     //                  .write
		.avmm_rcv_readdata    (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_readdata),  //                  .readdata
		.irq_space            (),                                                                //       (terminated)
		.irq_msg              ()                                                                 //       (terminated)
	);

	altera_avalon_mailbox #(
		.DWIDTH (32),
		.AWIDTH (2)
	) avalon_mailbox_out (
		.clk                  (clk_clk),                                                          //               clk.clk
		.rst_n                (~rst_controller_reset_out_reset),                                  //             rst_n.reset_n
		.avmm_snd_address     (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_address),     //   avmm_msg_sender.address
		.avmm_snd_writedata   (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_writedata),   //                  .writedata
		.avmm_snd_write       (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_write),       //                  .write
		.avmm_snd_read        (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_read),        //                  .read
		.avmm_snd_readdata    (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_readdata),    //                  .readdata
		.avmm_snd_waitrequest (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_waitrequest), //                  .waitrequest
		.avmm_rcv_address     (mailbox_out_address),                                              // avmm_msg_receiver.address
		.avmm_rcv_read        (mailbox_out_read),                                                 //                  .read
		.avmm_rcv_writedata   (mailbox_out_writedata),                                            //                  .writedata
		.avmm_rcv_write       (mailbox_out_write),                                                //                  .write
		.avmm_rcv_readdata    (mailbox_out_readdata),                                             //                  .readdata
		.irq_space            (),                                                                 //       (terminated)
		.irq_msg              ()                                                                  //       (terminated)
	);

	macci custom_instruction (
		.clk    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // nios_custom_instruction_slave.clk
		.clk_en (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.reset  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.n      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //                              .n
		.start  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.done   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.dataa  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //                              .dataa
		.datab  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                              .datab
		.result (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result)  //                              .result
	);

	multicore_system_core_0_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	multicore_system_core_1_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                                  clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                                reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                                     .reset_req
		.d_address                           (nios2_data_master_address),                           //                          data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (nios2_data_master_read),                              //                                     .read
		.d_readdata                          (nios2_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (nios2_data_master_write),                             //                                     .write
		.d_writedata                         (nios2_data_master_writedata),                         //                                     .writedata
		.d_burstcount                        (nios2_data_master_burstcount),                        //                                     .burstcount
		.d_readdatavalid                     (nios2_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                                     .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                                     .waitrequest
		.dtcm0_readdata                      (nios2_tightly_coupled_data_master_0_readdata),        //        tightly_coupled_data_master_0.readdata
		.dtcm0_address                       (nios2_tightly_coupled_data_master_0_address),         //                                     .address
		.dtcm0_read                          (nios2_tightly_coupled_data_master_0_read),            //                                     .read
		.dtcm0_clken                         (nios2_tightly_coupled_data_master_0_clken),           //                                     .clken
		.dtcm0_write                         (nios2_tightly_coupled_data_master_0_write),           //                                     .write
		.dtcm0_writedata                     (nios2_tightly_coupled_data_master_0_writedata),       //                                     .writedata
		.dtcm0_byteenable                    (nios2_tightly_coupled_data_master_0_byteenable),      //                                     .byteenable
		.itcm0_readdata                      (nios2_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (nios2_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (nios2_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (nios2_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.irq                                 (nios2_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                                     .writedata
		.A_ci_multi_done                     (nios2_custom_instruction_master_done),                //            custom_instruction_master.done
		.A_ci_multi_result                   (nios2_custom_instruction_master_multi_result),        //                                     .multi_result
		.A_ci_multi_a                        (nios2_custom_instruction_master_multi_a),             //                                     .multi_a
		.A_ci_multi_b                        (nios2_custom_instruction_master_multi_b),             //                                     .multi_b
		.A_ci_multi_c                        (nios2_custom_instruction_master_multi_c),             //                                     .multi_c
		.A_ci_multi_clk_en                   (nios2_custom_instruction_master_clk_en),              //                                     .clk_en
		.A_ci_multi_clock                    (nios2_custom_instruction_master_clk),                 //                                     .clk
		.A_ci_multi_reset                    (nios2_custom_instruction_master_reset),               //                                     .reset
		.A_ci_multi_reset_req                (nios2_custom_instruction_master_reset_req),           //                                     .reset_req
		.A_ci_multi_dataa                    (nios2_custom_instruction_master_multi_dataa),         //                                     .multi_dataa
		.A_ci_multi_datab                    (nios2_custom_instruction_master_multi_datab),         //                                     .multi_datab
		.A_ci_multi_n                        (nios2_custom_instruction_master_multi_n),             //                                     .multi_n
		.A_ci_multi_readra                   (nios2_custom_instruction_master_multi_readra),        //                                     .multi_readra
		.A_ci_multi_readrb                   (nios2_custom_instruction_master_multi_readrb),        //                                     .multi_readrb
		.A_ci_multi_start                    (nios2_custom_instruction_master_start),               //                                     .start
		.A_ci_multi_writerc                  (nios2_custom_instruction_master_multi_writerc)        //                                     .multi_writerc
	);

	multicore_system_core_3_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_1_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_1_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	multicore_system_core_3_rom rom (
		.address     (mm_interconnect_2_rom_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_rom_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_rom_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_rom_s1_write),      //       .write
		.readdata    (mm_interconnect_2_rom_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_rom_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_rom_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_rom_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_rom_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_rom_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_rom_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_rom_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_rom_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_rom_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                             //   clk1.clk
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	multicore_system_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                     //        ci_slave.result
		.ci_slave_multi_clk        (nios2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                     //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_n                (8'b00000000),                                                          //     (terminated)
		.ci_slave_readra           (1'b0),                                                                 //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                 //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                 //     (terminated)
		.ci_slave_a                (5'b00000),                                                             //     (terminated)
		.ci_slave_b                (5'b00000),                                                             //     (terminated)
		.ci_slave_c                (5'b00000),                                                             //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                 //     (terminated)
		.comb_ci_master_dataa      (),                                                                     //     (terminated)
		.comb_ci_master_datab      (),                                                                     //     (terminated)
		.comb_ci_master_n          (),                                                                     //     (terminated)
		.comb_ci_master_readra     (),                                                                     //     (terminated)
		.comb_ci_master_readrb     (),                                                                     //     (terminated)
		.comb_ci_master_writerc    (),                                                                     //     (terminated)
		.comb_ci_master_a          (),                                                                     //     (terminated)
		.comb_ci_master_b          (),                                                                     //     (terminated)
		.comb_ci_master_c          (),                                                                     //     (terminated)
		.comb_ci_master_ipending   (),                                                                     //     (terminated)
		.comb_ci_master_estatus    ()                                                                      //     (terminated)
	);

	multicore_system_core_0_nios2_custom_instruction_master_multi_xconnect nios2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (nios2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req ()                                                                          // (terminated)
	);

	multicore_system_core_0_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                  (clk_clk),                                                          //                           clock_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                   //   nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                      (nios2_data_master_address),                                        //                   nios2_data_master.address
		.nios2_data_master_waitrequest                  (nios2_data_master_waitrequest),                                    //                                    .waitrequest
		.nios2_data_master_burstcount                   (nios2_data_master_burstcount),                                     //                                    .burstcount
		.nios2_data_master_byteenable                   (nios2_data_master_byteenable),                                     //                                    .byteenable
		.nios2_data_master_read                         (nios2_data_master_read),                                           //                                    .read
		.nios2_data_master_readdata                     (nios2_data_master_readdata),                                       //                                    .readdata
		.nios2_data_master_readdatavalid                (nios2_data_master_readdatavalid),                                  //                                    .readdatavalid
		.nios2_data_master_write                        (nios2_data_master_write),                                          //                                    .write
		.nios2_data_master_writedata                    (nios2_data_master_writedata),                                      //                                    .writedata
		.nios2_data_master_debugaccess                  (nios2_data_master_debugaccess),                                    //                                    .debugaccess
		.nios2_instruction_master_address               (nios2_instruction_master_address),                                 //            nios2_instruction_master.address
		.nios2_instruction_master_waitrequest           (nios2_instruction_master_waitrequest),                             //                                    .waitrequest
		.nios2_instruction_master_read                  (nios2_instruction_master_read),                                    //                                    .read
		.nios2_instruction_master_readdata              (nios2_instruction_master_readdata),                                //                                    .readdata
		.avalon_data_bridge_s0_address                  (mm_interconnect_0_avalon_data_bridge_s0_address),                  //               avalon_data_bridge_s0.address
		.avalon_data_bridge_s0_write                    (mm_interconnect_0_avalon_data_bridge_s0_write),                    //                                    .write
		.avalon_data_bridge_s0_read                     (mm_interconnect_0_avalon_data_bridge_s0_read),                     //                                    .read
		.avalon_data_bridge_s0_readdata                 (mm_interconnect_0_avalon_data_bridge_s0_readdata),                 //                                    .readdata
		.avalon_data_bridge_s0_writedata                (mm_interconnect_0_avalon_data_bridge_s0_writedata),                //                                    .writedata
		.avalon_data_bridge_s0_burstcount               (mm_interconnect_0_avalon_data_bridge_s0_burstcount),               //                                    .burstcount
		.avalon_data_bridge_s0_byteenable               (mm_interconnect_0_avalon_data_bridge_s0_byteenable),               //                                    .byteenable
		.avalon_data_bridge_s0_readdatavalid            (mm_interconnect_0_avalon_data_bridge_s0_readdatavalid),            //                                    .readdatavalid
		.avalon_data_bridge_s0_waitrequest              (mm_interconnect_0_avalon_data_bridge_s0_waitrequest),              //                                    .waitrequest
		.avalon_data_bridge_s0_debugaccess              (mm_interconnect_0_avalon_data_bridge_s0_debugaccess),              //                                    .debugaccess
		.avalon_mailbox_in_avmm_msg_receiver_address    (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_address),    // avalon_mailbox_in_avmm_msg_receiver.address
		.avalon_mailbox_in_avmm_msg_receiver_write      (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_write),      //                                    .write
		.avalon_mailbox_in_avmm_msg_receiver_read       (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_read),       //                                    .read
		.avalon_mailbox_in_avmm_msg_receiver_readdata   (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_readdata),   //                                    .readdata
		.avalon_mailbox_in_avmm_msg_receiver_writedata  (mm_interconnect_0_avalon_mailbox_in_avmm_msg_receiver_writedata),  //                                    .writedata
		.avalon_mailbox_out_avmm_msg_sender_address     (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_address),     //  avalon_mailbox_out_avmm_msg_sender.address
		.avalon_mailbox_out_avmm_msg_sender_write       (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_write),       //                                    .write
		.avalon_mailbox_out_avmm_msg_sender_read        (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_read),        //                                    .read
		.avalon_mailbox_out_avmm_msg_sender_readdata    (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_readdata),    //                                    .readdata
		.avalon_mailbox_out_avmm_msg_sender_writedata   (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_writedata),   //                                    .writedata
		.avalon_mailbox_out_avmm_msg_sender_waitrequest (mm_interconnect_0_avalon_mailbox_out_avmm_msg_sender_waitrequest), //                                    .waitrequest
		.jtag_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_avalon_jtag_slave_address),                 //              jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_avalon_jtag_slave_write),                   //                                    .write
		.jtag_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_avalon_jtag_slave_read),                    //                                    .read
		.jtag_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                //                                    .readdata
		.jtag_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),               //                                    .writedata
		.jtag_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),             //                                    .waitrequest
		.jtag_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),              //                                    .chipselect
		.nios2_debug_mem_slave_address                  (mm_interconnect_0_nios2_debug_mem_slave_address),                  //               nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                    (mm_interconnect_0_nios2_debug_mem_slave_write),                    //                                    .write
		.nios2_debug_mem_slave_read                     (mm_interconnect_0_nios2_debug_mem_slave_read),                     //                                    .read
		.nios2_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_debug_mem_slave_readdata),                 //                                    .readdata
		.nios2_debug_mem_slave_writedata                (mm_interconnect_0_nios2_debug_mem_slave_writedata),                //                                    .writedata
		.nios2_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_debug_mem_slave_byteenable),               //                                    .byteenable
		.nios2_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),              //                                    .waitrequest
		.nios2_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),              //                                    .debugaccess
		.rom_s2_address                                 (mm_interconnect_0_rom_s2_address),                                 //                              rom_s2.address
		.rom_s2_write                                   (mm_interconnect_0_rom_s2_write),                                   //                                    .write
		.rom_s2_readdata                                (mm_interconnect_0_rom_s2_readdata),                                //                                    .readdata
		.rom_s2_writedata                               (mm_interconnect_0_rom_s2_writedata),                               //                                    .writedata
		.rom_s2_byteenable                              (mm_interconnect_0_rom_s2_byteenable),                              //                                    .byteenable
		.rom_s2_chipselect                              (mm_interconnect_0_rom_s2_chipselect),                              //                                    .chipselect
		.rom_s2_clken                                   (mm_interconnect_0_rom_s2_clken),                                   //                                    .clken
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                               //                            timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                                 //                                    .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                              //                                    .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                             //                                    .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect)                             //                                    .chipselect
	);

	multicore_system_core_0_mm_interconnect_1 mm_interconnect_1 (
		.clock_clk_clk                                  (clk_clk),                                        //                           clock_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                 //   nios2_reset_reset_bridge_in_reset.reset
		.nios2_tightly_coupled_data_master_0_address    (nios2_tightly_coupled_data_master_0_address),    // nios2_tightly_coupled_data_master_0.address
		.nios2_tightly_coupled_data_master_0_byteenable (nios2_tightly_coupled_data_master_0_byteenable), //                                    .byteenable
		.nios2_tightly_coupled_data_master_0_read       (nios2_tightly_coupled_data_master_0_read),       //                                    .read
		.nios2_tightly_coupled_data_master_0_readdata   (nios2_tightly_coupled_data_master_0_readdata),   //                                    .readdata
		.nios2_tightly_coupled_data_master_0_write      (nios2_tightly_coupled_data_master_0_write),      //                                    .write
		.nios2_tightly_coupled_data_master_0_writedata  (nios2_tightly_coupled_data_master_0_writedata),  //                                    .writedata
		.nios2_tightly_coupled_data_master_0_clken      (nios2_tightly_coupled_data_master_0_clken),      //                                    .clken
		.ram_s1_address                                 (mm_interconnect_1_ram_s1_address),               //                              ram_s1.address
		.ram_s1_write                                   (mm_interconnect_1_ram_s1_write),                 //                                    .write
		.ram_s1_readdata                                (mm_interconnect_1_ram_s1_readdata),              //                                    .readdata
		.ram_s1_writedata                               (mm_interconnect_1_ram_s1_writedata),             //                                    .writedata
		.ram_s1_byteenable                              (mm_interconnect_1_ram_s1_byteenable),            //                                    .byteenable
		.ram_s1_chipselect                              (mm_interconnect_1_ram_s1_chipselect),            //                                    .chipselect
		.ram_s1_clken                                   (mm_interconnect_1_ram_s1_clken)                  //                                    .clken
	);

	multicore_system_core_0_mm_interconnect_2 mm_interconnect_2 (
		.clock_clk_clk                                       (clk_clk),                                             //                                  clock_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                      //          nios2_reset_reset_bridge_in_reset.reset
		.nios2_tightly_coupled_instruction_master_0_address  (nios2_tightly_coupled_instruction_master_0_address),  // nios2_tightly_coupled_instruction_master_0.address
		.nios2_tightly_coupled_instruction_master_0_read     (nios2_tightly_coupled_instruction_master_0_read),     //                                           .read
		.nios2_tightly_coupled_instruction_master_0_readdata (nios2_tightly_coupled_instruction_master_0_readdata), //                                           .readdata
		.nios2_tightly_coupled_instruction_master_0_clken    (nios2_tightly_coupled_instruction_master_0_clken),    //                                           .clken
		.rom_s1_address                                      (mm_interconnect_2_rom_s1_address),                    //                                     rom_s1.address
		.rom_s1_write                                        (mm_interconnect_2_rom_s1_write),                      //                                           .write
		.rom_s1_readdata                                     (mm_interconnect_2_rom_s1_readdata),                   //                                           .readdata
		.rom_s1_writedata                                    (mm_interconnect_2_rom_s1_writedata),                  //                                           .writedata
		.rom_s1_byteenable                                   (mm_interconnect_2_rom_s1_byteenable),                 //                                           .byteenable
		.rom_s1_chipselect                                   (mm_interconnect_2_rom_s1_chipselect),                 //                                           .chipselect
		.rom_s1_clken                                        (mm_interconnect_2_rom_s1_clken)                       //                                           .clken
	);

	multicore_system_core_0_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
